module top;
  initial begin
    run_test("my_test");
  end
endmodule

/*
Concept
    -run_test() hands control to UVM
    -No manual instantiation
*/