package test_mode_pkg;
    typedef enum { SANITY, STRESS } test_mode_e;
endpackage