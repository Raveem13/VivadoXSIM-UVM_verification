interface my_if (input logic clk);
    logic rst;
    logic valid;
    logic [7:0] data;
endinterface //my_if 