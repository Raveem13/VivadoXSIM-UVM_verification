package test_mode_pkg;
    typedef enum { SANITY, STRESS, BURST } test_mode_e;
endpackage